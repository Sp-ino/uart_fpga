-- Copyright (c) 2023 Valerio Spinogatti
-- Licensed under Apache license

library ieee;
use ieee.std_logic_1164.all;


package common_pkg is

    constant byte_width_bit: integer := 8;
    constant word_width_byte: integer := 16;
    constant word_width_bit: integer := 128;

end common_pkg;